/vol/ece303/genus_tutorial/NangateOpenCellLibrary.lef
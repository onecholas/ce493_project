

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO eyeriss_top 
  PIN clk_i 
    ANTENNAPARTIALMETALAREA 9805.98 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 39533 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1439.76 LAYER metal3 ; 
    ANTENNAMAXAREACAR 50.3156 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 202.071 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.2058 LAYER via3 ;
    ANTENNAMAXCUTCAR 1.30681 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 15.3664 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 64.9936 LAYER metal4 ;
    ANTENNAGATEAREA 1612.04 LAYER metal4 ; 
    ANTENNAMAXAREACAR 50.3251 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 202.112 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0588 LAYER via4 ;
    ANTENNAMAXCUTCAR 1.30685 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.3132 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER metal5 ;
    ANTENNAGATEAREA 1612.2 LAYER metal5 ; 
    ANTENNAMAXAREACAR 50.326 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 202.115 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.30686 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 1.7444 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 7.056 LAYER metal6 ;
    ANTENNAGATEAREA 1612.27 LAYER metal6 ; 
    ANTENNAMAXAREACAR 50.327 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 202.119 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.30686 LAYER via6 ;
  END clk_i
  PIN rst_i 
    ANTENNAPARTIALMETALAREA 0.15295 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6118 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ; 
    ANTENNAMAXAREACAR 10.1733 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 40.5486 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.373333 LAYER via3 ;
  END rst_i
  PIN start_i 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END start_i
  PIN ifmap_wr_en_i 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.45742 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.7608 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END ifmap_wr_en_i
  PIN weight_wr_en_i 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_wr_en_i
  PIN ifmap_wr_addr_i[9] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.0439 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 48.5024 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_wr_addr_i[9]
  PIN ifmap_wr_addr_i[8] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_wr_addr_i[8]
  PIN ifmap_wr_addr_i[7] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 14 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 53.6244 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_wr_addr_i[7]
  PIN ifmap_wr_addr_i[6] 
    ANTENNAPARTIALMETALAREA 0.04655 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1862 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 14.9561 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 56.7073 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_wr_addr_i[6]
  PIN ifmap_wr_addr_i[5] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.45742 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.7608 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END ifmap_wr_addr_i[5]
  PIN ifmap_wr_addr_i[4] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ; 
    ANTENNAMAXAREACAR 10.4267 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 39.3638 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.373333 LAYER via3 ;
  END ifmap_wr_addr_i[4]
  PIN ifmap_wr_addr_i[3] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.522 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 50.4146 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_wr_addr_i[3]
  PIN ifmap_wr_addr_i[2] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4522 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 14.6488 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 56.2195 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_wr_addr_i[2]
  PIN ifmap_wr_addr_i[1] 
    ANTENNAPARTIALMETALAREA 0.04655 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1862 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 15.6049 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 59.1171 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_wr_addr_i[1]
  PIN ifmap_wr_addr_i[0] 
    ANTENNAPARTIALMETALAREA 0.07315 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.88 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 50.48 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.373333 LAYER via3 ;
  END ifmap_wr_addr_i[0]
  PIN ifmap_data_i[15] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.0976 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 41.2732 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[15]
  PIN ifmap_data_i[14] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[14]
  PIN ifmap_data_i[13] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3458 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 18.6098 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 72.4341 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[13]
  PIN ifmap_data_i[12] 
    ANTENNAPARTIALMETALAREA 0.05985 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2394 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.0098 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 49.6634 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[12]
  PIN ifmap_data_i[11] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[11]
  PIN ifmap_data_i[10] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.0976 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 41.2732 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[10]
  PIN ifmap_data_i[9] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[9]
  PIN ifmap_data_i[8] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3458 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.0537 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 46.2098 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[8]
  PIN ifmap_data_i[7] 
    ANTENNAPARTIALMETALAREA 0.04655 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1862 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 15.4341 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 58.6195 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[7]
  PIN ifmap_data_i[6] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[6]
  PIN ifmap_data_i[5] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.0976 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 41.2732 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[5]
  PIN ifmap_data_i[4] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[4]
  PIN ifmap_data_i[3] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3458 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.0537 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 46.2098 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[3]
  PIN ifmap_data_i[2] 
    ANTENNAPARTIALMETALAREA 0.07315 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.0098 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 49.8488 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[2]
  PIN ifmap_data_i[1] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[1]
  PIN ifmap_data_i[0] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.0976 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 41.2732 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END ifmap_data_i[0]
  PIN weight_data_i[15] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.0976 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 41.2732 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[15]
  PIN weight_data_i[14] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[14]
  PIN weight_data_i[13] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3458 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.0537 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 46.2098 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[13]
  PIN weight_data_i[12] 
    ANTENNAPARTIALMETALAREA 0.07315 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.4878 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 51.761 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[12]
  PIN weight_data_i[11] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.9659 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 54.0439 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[11]
  PIN weight_data_i[10] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.0976 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 41.2732 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[10]
  PIN weight_data_i[9] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[9]
  PIN weight_data_i[8] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.0537 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 46.3951 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[8]
  PIN weight_data_i[7] 
    ANTENNAPARTIALMETALAREA 0.04655 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1862 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.4878 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 51.3902 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[7]
  PIN weight_data_i[6] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3458 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.9659 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 53.8585 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[6]
  PIN weight_data_i[5] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.0976 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 41.2732 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[5]
  PIN weight_data_i[4] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[4]
  PIN weight_data_i[3] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3458 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.0537 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 46.2098 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[3]
  PIN weight_data_i[2] 
    ANTENNAPARTIALMETALAREA 0.04655 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1862 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.0098 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 49.478 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[2]
  PIN weight_data_i[1] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[1]
  PIN weight_data_i[0] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.0976 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 41.2732 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_data_i[0]
  PIN weight_wr_addr_i[4] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.0976 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 41.2732 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_wr_addr_i[4]
  PIN weight_wr_addr_i[3] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5756 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 43.1854 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_wr_addr_i[3]
  PIN weight_wr_addr_i[2] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.0537 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 46.3951 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_wr_addr_i[2]
  PIN weight_wr_addr_i[1] 
    ANTENNAPARTIALMETALAREA 0.05985 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2394 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.4878 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 51.5756 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_wr_addr_i[1]
  PIN weight_wr_addr_i[0] 
    ANTENNAPARTIALMETALAREA 0.00665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0266 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.522 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 50.4146 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.478049 LAYER via3 ;
  END weight_wr_addr_i[0]
  PIN psum_rd_en_i[0] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.418 LAYER metal3 ; 
    ANTENNAMAXAREACAR 1.25263 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 4.88732 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.023445 LAYER via3 ;
  END psum_rd_en_i[0]
  PIN psum_rd_en_i[1] 
    ANTENNAPARTIALMETALAREA 0.24605 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9842 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.836 LAYER metal3 ; 
    ANTENNAMAXAREACAR 1.32679 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 4.4756 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.0117225 LAYER via3 ;
  END psum_rd_en_i[1]
  PIN psum_rd_en_i[2] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.672 LAYER metal3 ; 
    ANTENNAMAXAREACAR 0.881699 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 3.35574 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.00586124 LAYER via3 ;
  END psum_rd_en_i[2]
  PIN psum_rd_en_i[3] 
    ANTENNAPARTIALMETALAREA 0.28595 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1438 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.836 LAYER metal3 ; 
    ANTENNAMAXAREACAR 1.23433 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 4.1116 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.0117225 LAYER via3 ;
  END psum_rd_en_i[3]
  PIN psum_rd_en_i[4] 
    ANTENNAPARTIALMETALAREA 0.25935 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0374 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.836 LAYER metal3 ; 
    ANTENNAMAXAREACAR 2.05197 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 7.37739 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.0117225 LAYER via3 ;
  END psum_rd_en_i[4]
  PIN psum_rd_en_i[5] 
    ANTENNAPARTIALMETALAREA 0.33565 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3426 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.836 LAYER metal3 ; 
    ANTENNAMAXAREACAR 1.76394 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 6.22524 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.0117225 LAYER via3 ;
  END psum_rd_en_i[5]
  PIN psum_empty_o[0] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1372 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5684 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.3524 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.1155 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 4.4884 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 18.032 LAYER metal6 ;
  END psum_empty_o[0]
  PIN psum_empty_o[1] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1372 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5684 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.3516 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.4848 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.202125 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 21.8148 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 87.3376 LAYER metal6 ;
  END psum_empty_o[1]
  PIN psum_empty_o[2] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.49 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9796 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.4308 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8016 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.202125 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 16.4444 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 65.856 LAYER metal6 ;
  END psum_empty_o[2]
  PIN psum_empty_o[3] 
    ANTENNAPARTIALMETALAREA 0.10955 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4069 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2058 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8428 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.274 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1744 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 12.9948 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 52.0576 LAYER metal6 ;
  END psum_empty_o[3]
  PIN psum_empty_o[4] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.784 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.1463 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 34.2804 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 137.2 LAYER metal6 ;
  END psum_empty_o[4]
  PIN psum_empty_o[5] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.202125 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 33.6728 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 134.848 LAYER metal6 ;
  END psum_empty_o[5]
  PIN psum_o\[5\][15] 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.6608 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6628 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.3524 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4292 LAYER metal3 ;
  END psum_o\[5\][15]
  PIN psum_o\[5\][14] 
    ANTENNAPARTIALMETALAREA 0.28595 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0621 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.301 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2236 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.1095 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4576 LAYER metal3 ;
  END psum_o\[5\][14]
  PIN psum_o\[5\][13] 
    ANTENNAPARTIALMETALAREA 0.17955 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6669 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3255 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3412 LAYER metal3 ;
  END psum_o\[5\][13]
  PIN psum_o\[5\][12] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4199 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3892 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5764 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2226 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.91 LAYER metal3 ;
  END psum_o\[5\][12]
  PIN psum_o\[5\][11] 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4693 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3332 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3524 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.2859 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1632 LAYER metal3 ;
  END psum_o\[5\][11]
  PIN psum_o\[5\][10] 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4693 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4018 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6268 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.89275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.6102 LAYER metal3 ;
  END psum_o\[5\][10]
  PIN psum_o\[5\][9] 
    ANTENNAPARTIALMETALAREA 0.40565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5067 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3724 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5092 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5278 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1308 LAYER metal3 ;
  END psum_o\[5\][9]
  PIN psum_o\[5\][8] 
    ANTENNAPARTIALMETALAREA 0.62475 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3205 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.049 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2156 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.5526 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.23 LAYER metal3 ;
  END psum_o\[5\][8]
  PIN psum_o\[5\][7] 
    ANTENNAPARTIALMETALAREA 0.30205 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1219 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3486 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.414 LAYER metal3 ;
  END psum_o\[5\][7]
  PIN psum_o\[5\][6] 
    ANTENNAPARTIALMETALAREA 0.31885 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1843 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2023 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8288 LAYER metal3 ;
  END psum_o\[5\][6]
  PIN psum_o\[5\][5] 
    ANTENNAPARTIALMETALAREA 0.28595 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0621 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0203 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1008 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.086625 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 1.6072 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5072 LAYER metal4 ;
  END psum_o\[5\][5]
  PIN psum_o\[5\][4] 
    ANTENNAPARTIALMETALAREA 1.09725 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0755 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.1364 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5848 LAYER metal3 ;
  END psum_o\[5\][4]
  PIN psum_o\[5\][3] 
    ANTENNAPARTIALMETALAREA 0.33915 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2597 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2681 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.092 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2289 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9352 LAYER metal3 ;
  END psum_o\[5\][3]
  PIN psum_o\[5\][2] 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4693 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2548 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.004 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0356 LAYER metal3 ;
  END psum_o\[5\][2]
  PIN psum_o\[5\][1] 
    ANTENNAPARTIALMETALAREA 0.21945 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8151 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 3.0436 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.194 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.7538 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.0348 LAYER metal3 ;
  END psum_o\[5\][1]
  PIN psum_o\[5\][0] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.6468 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6068 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.4116 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 7.7028 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 30.8896 LAYER metal6 ;
  END psum_o\[5\][0]
  PIN psum_o\[4\][15] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4116 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 8.2908 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 33.2416 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.1155 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.1364 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.624 LAYER metal6 ;
  END psum_o\[4\][15]
  PIN psum_o\[4\][14] 
    ANTENNAPARTIALMETALAREA 0.18585 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6903 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0329 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1512 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 3.6057 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.4424 LAYER metal3 ;
  END psum_o\[4\][14]
  PIN psum_o\[4\][13] 
    ANTENNAPARTIALMETALAREA 0.20895 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7761 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 3.3026 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.2496 LAYER metal3 ;
  END psum_o\[4\][13]
  PIN psum_o\[4\][12] 
    ANTENNAPARTIALMETALAREA 0.41195 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5301 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 3.3418 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3868 LAYER metal3 ;
  END psum_o\[4\][12]
  PIN psum_o\[4\][11] 
    ANTENNAPARTIALMETALAREA 0.13965 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5187 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1764 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3521 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4476 LAYER metal3 ;
  END psum_o\[4\][11]
  PIN psum_o\[4\][10] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4872 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9684 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4151 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER metal3 ;
  END psum_o\[4\][10]
  PIN psum_o\[4\][9] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3211 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2156 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0238 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1148 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.9604 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.92 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.7636 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 11.1328 LAYER metal6 ;
  END psum_o\[4\][9]
  PIN psum_o\[4\][8] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4116 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 2.9596 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 11.9168 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.1155 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.626 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 14.5824 LAYER metal6 ;
  END psum_o\[4\][8]
  PIN psum_o\[4\][7] 
    ANTENNAPARTIALMETALAREA 0.20615 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7657 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.812 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.086625 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 2.4108 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.7216 LAYER metal4 ;
  END psum_o\[4\][7]
  PIN psum_o\[4\][6] 
    ANTENNAPARTIALMETALAREA 0.27265 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0127 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3332 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.329 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3356 LAYER metal3 ;
  END psum_o\[4\][6]
  PIN psum_o\[4\][5] 
    ANTENNAPARTIALMETALAREA 0.35245 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3091 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8036 LAYER metal3 ;
  END psum_o\[4\][5]
  PIN psum_o\[4\][4] 
    ANTENNAPARTIALMETALAREA 0.17255 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6409 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2548 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4683 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8928 LAYER metal3 ;
  END psum_o\[4\][4]
  PIN psum_o\[4\][3] 
    ANTENNAPARTIALMETALAREA 0.10955 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4069 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3598 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1162 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4844 LAYER metal3 ;
  END psum_o\[4\][3]
  PIN psum_o\[4\][2] 
    ANTENNAPARTIALMETALAREA 0.26565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9867 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.8204 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3012 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2093 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8568 LAYER metal3 ;
  END psum_o\[4\][2]
  PIN psum_o\[4\][1] 
    ANTENNAPARTIALMETALAREA 0.17955 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6669 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.61055 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.4618 LAYER metal3 ;
  END psum_o\[4\][1]
  PIN psum_o\[4\][0] 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4693 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.6758 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7228 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1029 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4312 LAYER metal3 ;
  END psum_o\[4\][0]
  PIN psum_o\[3\][15] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4199 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3402 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3804 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2226 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.91 LAYER metal3 ;
  END psum_o\[3\][15]
  PIN psum_o\[3\][14] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4199 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.6342 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5564 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2359 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9632 LAYER metal3 ;
  END psum_o\[3\][14]
  PIN psum_o\[3\][13] 
    ANTENNAPARTIALMETALAREA 0.13615 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5057 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.086625 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 0.9513 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8248 LAYER metal2 ;
  END psum_o\[3\][13]
  PIN psum_o\[3\][12] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3211 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.497 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0076 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0238 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1148 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.0188 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1536 LAYER metal6 ;
  END psum_o\[3\][12]
  PIN psum_o\[3\][11] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3211 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5236 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.114 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.5253 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1208 LAYER metal3 ;
  END psum_o\[3\][11]
  PIN psum_o\[3\][10] 
    ANTENNAPARTIALMETALAREA 0.18585 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6903 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4053 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6604 LAYER metal3 ;
  END psum_o\[3\][10]
  PIN psum_o\[3\][9] 
    ANTENNAPARTIALMETALAREA 0.33845 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2571 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.086625 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 0.2422 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9884 LAYER metal2 ;
  END psum_o\[3\][9]
  PIN psum_o\[3\][8] 
    ANTENNAPARTIALMETALAREA 0.15925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5915 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3332 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4753 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9208 LAYER metal3 ;
  END psum_o\[3\][8]
  PIN psum_o\[3\][7] 
    ANTENNAPARTIALMETALAREA 0.17955 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6669 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1561 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER metal3 ;
  END psum_o\[3\][7]
  PIN psum_o\[3\][6] 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4693 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.1368 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5668 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4487 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8144 LAYER metal3 ;
  END psum_o\[3\][6]
  PIN psum_o\[3\][5] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3211 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4774 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9292 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4284 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7332 LAYER metal3 ;
  END psum_o\[3\][5]
  PIN psum_o\[3\][4] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.7126 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.784 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.5476 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 14.2688 LAYER metal6 ;
  END psum_o\[3\][4]
  PIN psum_o\[3\][3] 
    ANTENNAPARTIALMETALAREA 0.24605 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9139 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.9282 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7324 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1029 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4312 LAYER metal3 ;
  END psum_o\[3\][3]
  PIN psum_o\[3\][2] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4199 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0168 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0868 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1.7052 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8992 LAYER metal6 ;
  END psum_o\[3\][2]
  PIN psum_o\[3\][1] 
    ANTENNAPARTIALMETALAREA 0.20615 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7657 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1827 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7504 LAYER metal3 ;
  END psum_o\[3\][1]
  PIN psum_o\[3\][0] 
    ANTENNAPARTIALMETALAREA 0.26565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9867 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5754 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3212 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2891 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.176 LAYER metal3 ;
  END psum_o\[3\][0]
  PIN psum_o\[2\][15] 
    ANTENNAPARTIALMETALAREA 0.24885 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9243 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.9702 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9004 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3423 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3888 LAYER metal3 ;
  END psum_o\[2\][15]
  PIN psum_o\[2\][14] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.504 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0356 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2548 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0976 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.4484 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 25.872 LAYER metal6 ;
  END psum_o\[2\][14]
  PIN psum_o\[2\][13] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4199 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.086625 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 1.4308 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7428 LAYER metal2 ;
  END psum_o\[2\][13]
  PIN psum_o\[2\][12] 
    ANTENNAPARTIALMETALAREA 0.19285 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7163 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.2114 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8652 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.086625 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 1.3328 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4096 LAYER metal4 ;
  END psum_o\[2\][12]
  PIN psum_o\[2\][11] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4382 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7724 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.9569 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8472 LAYER metal3 ;
  END psum_o\[2\][11]
  PIN psum_o\[2\][10] 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4693 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1274 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5292 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1561 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER metal3 ;
  END psum_o\[2\][10]
  PIN psum_o\[2\][9] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4199 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1764 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4018 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6268 LAYER metal3 ;
  END psum_o\[2\][9]
  PIN psum_o\[2\][8] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4018 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6268 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.3552 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4404 LAYER metal3 ;
  END psum_o\[2\][8]
  PIN psum_o\[2\][7] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4746 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5145 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0776 LAYER metal3 ;
  END psum_o\[2\][7]
  PIN psum_o\[2\][6] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4199 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3794 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5372 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4613 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8648 LAYER metal3 ;
  END psum_o\[2\][6]
  PIN psum_o\[2\][5] 
    ANTENNAPARTIALMETALAREA 0.09625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3575 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.6048 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4388 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.3766 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.526 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.7252 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9792 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1.9012 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6832 LAYER metal6 ;
  END psum_o\[2\][5]
  PIN psum_o\[2\][4] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1176 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.49 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 7.7812 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 31.2032 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 0.9212 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7632 LAYER metal6 ;
  END psum_o\[2\][4]
  PIN psum_o\[2\][3] 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4693 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3626 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.47 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.1531 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.632 LAYER metal3 ;
  END psum_o\[2\][3]
  PIN psum_o\[2\][2] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3211 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5684 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2932 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1295 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5376 LAYER metal3 ;
  END psum_o\[2\][2]
  PIN psum_o\[2\][1] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3211 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5488 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2148 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0238 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1148 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1.862 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5264 LAYER metal6 ;
  END psum_o\[2\][1]
  PIN psum_o\[2\][0] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.086625 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 0.7287 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9344 LAYER metal2 ;
  END psum_o\[2\][0]
  PIN psum_o\[1\][15] 
    ANTENNAPARTIALMETALAREA 0.24605 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9139 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3304 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3412 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.5472 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.228 LAYER metal3 ;
  END psum_o\[1\][15]
  PIN psum_o\[1\][14] 
    ANTENNAPARTIALMETALAREA 0.20615 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7657 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3689 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4952 LAYER metal3 ;
  END psum_o\[1\][14]
  PIN psum_o\[1\][13] 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4693 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3332 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4151 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER metal3 ;
  END psum_o\[1\][13]
  PIN psum_o\[1\][12] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3211 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.086625 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 1.799 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2156 LAYER metal2 ;
  END psum_o\[1\][12]
  PIN psum_o\[1\][11] 
    ANTENNAPARTIALMETALAREA 0.11935 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4433 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.086625 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 0.9219 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7072 LAYER metal2 ;
  END psum_o\[1\][11]
  PIN psum_o\[1\][10] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4199 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4998 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0188 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1694 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6972 LAYER metal3 ;
  END psum_o\[1\][10]
  PIN psum_o\[1\][9] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1568 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6468 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.49 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0384 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.8812 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 11.6032 LAYER metal6 ;
  END psum_o\[1\][9]
  PIN psum_o\[1\][8] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4116 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.4692 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.9552 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.5676 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3488 LAYER metal6 ;
  END psum_o\[1\][8]
  PIN psum_o\[1\][7] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4199 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1764 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0168 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0868 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.784 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.4892 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0352 LAYER metal6 ;
  END psum_o\[1\][7]
  PIN psum_o\[1\][6] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4199 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.448 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8116 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3822 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5484 LAYER metal3 ;
  END psum_o\[1\][6]
  PIN psum_o\[1\][5] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3332 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 2.3617 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.7406 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.982 LAYER metal3 ;
  END psum_o\[1\][5]
  PIN psum_o\[1\][4] 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4693 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0686 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.294 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3689 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4952 LAYER metal3 ;
  END psum_o\[1\][4]
  PIN psum_o\[1\][3] 
    ANTENNAPARTIALMETALAREA 0.39235 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4573 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3619 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4672 LAYER metal3 ;
  END psum_o\[1\][3]
  PIN psum_o\[1\][2] 
    ANTENNAPARTIALMETALAREA 0.17255 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6409 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.329 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3356 LAYER metal3 ;
  END psum_o\[1\][2]
  PIN psum_o\[1\][1] 
    ANTENNAPARTIALMETALAREA 0.36855 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3689 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.9931 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.0116 LAYER metal3 ;
  END psum_o\[1\][1]
  PIN psum_o\[1\][0] 
    ANTENNAPARTIALMETALAREA 0.23905 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8879 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4116 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.666 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.8141 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.276 LAYER metal3 ;
  END psum_o\[1\][0]
  PIN psum_o\[0\][15] 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.086625 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 0.9254 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7212 LAYER metal2 ;
  END psum_o\[0\][15]
  PIN psum_o\[0\][14] 
    ANTENNAPARTIALMETALAREA 0.24605 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9139 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.086625 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 1.2264 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9252 LAYER metal2 ;
  END psum_o\[0\][14]
  PIN psum_o\[0\][13] 
    ANTENNAPARTIALMETALAREA 0.21945 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8151 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.086625 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 0.147 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6076 LAYER metal2 ;
  END psum_o\[0\][13]
  PIN psum_o\[0\][12] 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4693 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3234 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3132 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5215 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1056 LAYER metal3 ;
  END psum_o\[0\][12]
  PIN psum_o\[0\][11] 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2191 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.896 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.6111 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.464 LAYER metal3 ;
  END psum_o\[0\][11]
  PIN psum_o\[0\][10] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2744 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1172 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.3524 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.9004 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 15.68 LAYER metal6 ;
  END psum_o\[0\][10]
  PIN psum_o\[0\][9] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5894 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3772 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.8228 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3696 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 1.1704 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.4684 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.952 LAYER metal6 ;
  END psum_o\[0\][9]
  PIN psum_o\[0\][8] 
    ANTENNAPARTIALMETALAREA 0.22575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8385 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.2177 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8904 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.086625 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 2.254 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.0944 LAYER metal4 ;
  END psum_o\[0\][8]
  PIN psum_o\[0\][7] 
    ANTENNAPARTIALMETALAREA 0.20895 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7761 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.086625 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 0.5859 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3632 LAYER metal2 ;
  END psum_o\[0\][7]
  PIN psum_o\[0\][6] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4199 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.49 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9796 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2359 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9632 LAYER metal3 ;
  END psum_o\[0\][6]
  PIN psum_o\[0\][5] 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3211 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.35 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4196 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.5225 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1096 LAYER metal3 ;
  END psum_o\[0\][5]
  PIN psum_o\[0\][4] 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3705 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.6671 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.688 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0105 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.8428 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4496 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.086625 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.0972 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.4672 LAYER metal6 ;
  END psum_o\[0\][4]
  PIN psum_o\[0\][3] 
    ANTENNAPARTIALMETALAREA 0.13965 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5187 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2758 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1228 LAYER metal3 ;
  END psum_o\[0\][3]
  PIN psum_o\[0\][2] 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4693 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1372 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.2387 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9744 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.086625 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 2.5676 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3488 LAYER metal4 ;
  END psum_o\[0\][2]
  PIN psum_o\[0\][1] 
    ANTENNAPARTIALMETALAREA 0.16625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6175 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.02205 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1078 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.7038 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8348 LAYER metal3 ;
  END psum_o\[0\][1]
  PIN psum_o\[0\][0] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4199 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.7098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.086625 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.8008 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2228 LAYER metal3 ;
  END psum_o\[0\][0]
END eyeriss_top

END LIBRARY
